LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
ENTITY bcd1 IS
PORT
(Q:IN STD_LOGIC_VECTOR(3 downto 0);
 P1,P2:BUFFER STD_LOGIC_VECTOR(3 downto 0);
 C0:OUT STD_LOGIC_VECTOR(7 downto 0);
 C1:OUT STD_LOGIC_VECTOR(7 downto 0)
 );
END bcd1;

ARCHITECTURE behave OF bcd1 IS
BEGIN
process(Q)
BEGIN
CASE Q IS
  WHEN "0000"=>P1<="0000";P2<="0000";
  WHEN "0001"=>P1<="0001";P2<="0000";
  WHEN "0010"=>P1<="0010";P2<="0000";
  WHEN "0011"=>P1<="0011";P2<="0000";
  WHEN "0100"=>P1<="0100";P2<="0000";
  WHEN "0101"=>P1<="0101";P2<="0000";
  WHEN "0110"=>P1<="0110";P2<="0000";
  WHEN "0111"=>P1<="0111";P2<="0000";
  WHEN "1000"=>P1<="1000";P2<="0000";
  WHEN "1001"=>P1<="1001";P2<="0000";
  WHEN "1010"=>P1<="0000";P2<="0001";
  WHEN "1011"=>P1<="0001";P2<="0001"; 
  WHEN "1100"=>P1<="0010";P2<="0001"; 
  WHEN "1101"=>P1<="0011";P2<="0001";
  WHEN "1110"=>P1<="0100";P2<="0001";
  WHEN "1111"=>P1<="0101";P2<="0001";
  WHEN others=>null;
END CASE;
CASE P1 IS
 WHEN "0000"=>C1<="11000000";     
 WHEN "0001"=>C1<="11111001";
 WHEN "0010"=>C1<="10100100";
 WHEN "0011"=>C1<="10110000";
 WHEN "0100"=>C1<="10011001";
 WHEN "0101"=>C1<="10010010";
 WHEN "0110"=>C1<="10000010";
 WHEN "0111"=>C1<="11111000";
 WHEN "1000"=>C1<="10000000";
 WHEN "1001"=>C1<="10010000";
 WHEN others=>null;
END CASE; 
CASE P2 IS
 WHEN "0000"=>C0<="11000000";     
 WHEN "0001"=>C0<="11111001";
 WHEN "0010"=>C0<="10100100";
 WHEN "0011"=>C0<="10110000";
 WHEN "0100"=>C0<="10011001";
 WHEN "0101"=>C0<="10010010";
 WHEN "0110"=>C0<="10000010";
 WHEN "0111"=>C0<="11111000";
 WHEN "1000"=>C0<="10000000";
 WHEN "1001"=>C0<="10010000";
 WHEN others=>null;
END CASE; 

end process;
END behave;